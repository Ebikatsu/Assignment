module sevenseg(input logic [3:0]data,
		output logic [6:0]segments);
	always_comb
	case(data)
		4'h0: segments = 7'b111_1110;
		4'h1: segments = 7'b011_0000;
		4'h2: segments = 7'b110_1101;
		4'h3: segments = 7'b111_1001;
		4'h4: segments = 7'b011_0011;
		4'h5: segments = 7'b101_1011;
		4'h6: segments = 7'b101_1111;
		4'h7: segments = 7'b111_0000;
		4'h8: segments = 7'b111_1111;
		4'h9: segments = 7'b111_0011;
		4'ha: segments = 7'b111_0111;
		4'hb: segments = 7'b001_1111;
		4'hc: segments = 7'b100_1110;
		4'hd: segments = 7'b011_1101;
		4'he: segments = 7'b100_1111;
		4'hf: segments = 7'b100_0111;
	endcase
endmodule
