module testbench();
	logic	clk50;
	logic	clk1;
	clkgen1m clkgen1m(clk50,clk1);
	initial begin
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
		clk50=0;#10;
		clk50=1;#10;
	end
endmodule
